// program counter
// supports both relative and absolute jumps
// use either or both, as desired
module PC #(parameter D=10)(
  input reset,					// synchronous reset
        clk,
        // reljump_en,             // rel. jump enable
        absjump_en,				// abs. jump enable
        jmp_en,
  input       [D-1:0] target,	// how far/where to jump
  input       [D-1:0] absaddress,
  output logic[D-1:0] prog_ctr
);


  always_ff @(posedge clk) begin
    if(reset)
	    prog_ctr <= 'b0;
    // else if(reljump_en)
      // prog_ctr <= prog_ctr + target;
    else if(jmp_en && absjump_en)
	    prog_ctr <= absaddress;
    else if(jmp_en)
      prog_ctr <= prog_ctr + target;
    else
      prog_ctr <= prog_ctr + 'b1;
  end

endmodule